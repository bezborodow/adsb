library ieee;                        
use ieee.std_logic_1164.all;         
use ieee.numeric_std.all;            

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package adsb_pkg is
    constant DEFAULT_SAMPLES_PER_SYMBOL    : integer := 10;
    constant DEFAULT_BUFFER_SYMBOL_LENGTH  : integer := 16;
    constant DEFAULT_IQ_WIDTH              : integer := 12;
end package adsb_pkg;

package body adsb_pkg is
end package body adsb_pkg;
